library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
 
entity hazard_detection_unit is
	 Port ( 

	 );
	 
	 
end alu;
 
architecture arch of hazard_detection_unit is

	
begin
	process(all) begin
		
	end process;
end architecture;